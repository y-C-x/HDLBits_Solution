module top_module (
    input a,
    input b,
    input c,
    input d,
    output q );//

    assign q = b & (d | c) | a & (c | d); // Fix me

endmodule
